���.      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.2.2�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby_wsp��wzrost��leki�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh&hNhJ�
hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h4�f8�����R�(KhKNNNJ����J����K t�b�C              �?�t�bhOh(�scalar���hJC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hK�
node_count�K�nodes�h*h-K ��h/��R�(KK��h4�V56�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h{h4�i8�����R�(KhKNNNJ����J����K t�bK ��h|h�K��h}h�K��h~h[K��hh[K ��h�h�K(��h�h[K0��uK8KKt�b�Bh                            �@@�q�q�?             H@                           �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?                            @>A�F<�?             C@                          ph@     ��?             @@������������������������       �                     =@������������������������       �                     @	       
                   �P@�q�q�?             @������������������������       �z�G�z�?             @������������������������       �                     �?�t�b�values�h*h-K ��h/��R�(KKKK��h[�C�      @@      0@      �?      "@              "@      �?              ?@      @      =@      @      =@                      @       @      @      �?      @      �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ/��hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�BH                            pg@r�q��?!             H@                          �E@X�Cc�?             <@                         �uf@X�Cc�?             ,@������������������������       �؇���X�?             @������������������������       �և���X�?             @                            @@4և���?             ,@������������������������       �        	             (@������������������������       �      �?              @	                           �?z�G�z�?             4@
                          �C@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @                          �0@      �?
             0@������������������������       �                     �?������������������������       ���S�ۿ?	             .@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      6@      :@      2@      $@      @      "@      �?      @      @      @      *@      �?      (@              �?      �?      @      0@       @       @              �?       @      �?       @      ,@      �?              �?      ,@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJu�7hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�Bh                            �E@�q���?             H@                           @�X�<ݺ?
             2@������������������������       �                     0@                          �g@      �?              @������������������������       �                     �?������������������������       �                     �?       
                   �g@������?             >@       	                  �%g@�8��8��?             8@������������������������       �        
             0@������������������������       �      �?              @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      7@      9@      �?      1@              0@      �?      �?              �?      �?              6@       @      6@       @      0@              @       @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ��!XhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                              �?r�q��?             H@������������������������       �                     &@                          �h@�Gi����?            �B@                          �@@�g�y��?             ?@������������������������       �8�Z$���?             *@������������������������       ��E��ӭ�?             2@������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�Cp      :@      6@      &@              .@      6@      .@      0@       @      &@      *@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJC�NhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrK	hsh*h-K ��h/��R�(KK	��hz�B�                             @�q�q�?#             H@                          �g@�eP*L��?!             F@                            @:ɨ��?            �@@������������������������       ��J�4�?             9@������������������������       �      �?              @                           @�C��2(�?
             &@������������������������       �        	             $@������������������������       �                     �?������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK	KK��h[�C�      <@      4@      8@      4@      7@      $@      5@      @       @      @      �?      $@              $@      �?              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�R�[hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�Bh                            �E@      �?             H@                          pg@�X����?             6@                           @���|���?             &@������������������������       �X�<ݚ�?             "@������������������������       �                      @������������������������       �                     &@       
                   �g@ȵHPS!�?             :@       	                     @ �q�q�?             8@������������������������       �                     3@������������������������       �z�G�z�?             @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      >@      2@      @      .@      @      @      @      @       @                      &@      7@      @      7@      �?      3@              @      �?               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�v}hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrK	hsh*h-K ��h/��R�(KK	��hz�B�                            �@@     ��?             H@������������������������       �                     *@                          �E@4�2%ޑ�?            �A@                          �g@      �?              @������������������������       �z�G�z�?             @������������������������       �                     @                           R@PN��T'�?             ;@������������������������       ����}<S�?             7@������������������������       �      �?             @�t�bh�h*h-K ��h/��R�(KK	KK��h[�C�      ;@      5@              *@      ;@       @      @      @      �?      @      @              7@      @      5@       @       @       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJg}�XhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrK	hsh*h-K ��h/��R�(KK	��hz�B�                            �h@      �?             H@                            @����X�?             E@                         ��f@4�2%ޑ�?            �A@������������������������       ��KM�]�?             3@������������������������       �      �?	             0@                           @և���X�?             @������������������������       �      �?             @������������������������       �                     @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK	KK��h[�C�      >@      2@      >@      (@      ;@       @      1@       @      $@      @      @      @      @      �?              @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ	�tlhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�Bh                              �?     ��?             H@                          �g@؇���X�?             ,@������������������������       �                     (@������������������������       �                      @                           @�������?             A@                           0@j���� �?             1@������������������������       �                      @������������������������       ��q�q�?             .@	       
                   �d@�t����?
             1@������������������������       �                     �?������������������������       �      �?	             0@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      5@      ;@      (@       @      (@                       @      "@      9@      @      $@       @              @      $@       @      .@      �?              �?      .@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�ޡhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                           y�E@�q���?             H@                           @������?             >@                          �g@��s����?             5@������������������������       ����|���?             &@������������������������       �                     $@                           �?X�<ݚ�?             "@������������������������       �����X�?             @������������������������       �                      @	       
                    @�X�<ݺ?             2@������������������������       �                     (@                           �?r�q��?             @������������������������       �      �?              @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      9@      7@       @      6@      @      1@      @      @              $@      @      @       @      @       @              1@      �?      (@              @      �?      �?      �?      @        �t�bubhhubehhub.